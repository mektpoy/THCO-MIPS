library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Controller is
    Port 
    ( 
		instrId : in STD_LOGIC_VECTOR (4 downto 0);
		stay : in STD_LOGIC;
		aluOp : out STD_LOGIC_VECTOR (2 downto 0);
		BMuxOp : out STD_LOGIC;
		jumpType : out STD_LOGIC_VECTOR (2 downto 0);
		resultSrc : out STD_LOGIC;
		memoryMode : out STD_LOGIC_VECTOR (1 downto 0);
		aluResultSrc : out STD_LOGIC_VECTOR (1 downto 0);
		regWrite : out STD_LOGIC;
		memoryRead : out STD_LOGIC
	);
end Controller;

architecture Behavioral of Controller is
begin
	process (instrId, stay)
	begin
		if (stay = '1') then
			aluOp <= "111";
			BMuxOp <= '0';
			jumpType <= "000";
			resultSrc <= '1';
			memoryMode <= "00";
			aluResultSrc <= "10";
			regWrite <= '0';
			memoryRead <= '0';
		else
			case instrId is
				when "00001" => -- ADDIU
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "00010" => -- ADDIU3
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "00011" => -- ADDSP3
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "00100" => -- ADDSP
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "00101" => -- ADDU
					aluOp <= "000";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "00110" => -- AND
					aluOp <= "010";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "00111" => -- B
					aluOp <= "111";
					BMuxOp <= '1';
					jumpType <= "001";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '0';
					memoryRead <= '0';
				when "01000" => -- BEQZ
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "010";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '0';
					memoryRead <= '0';
				when "01001" => -- BNEZ
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "011";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '0';
					memoryRead <= '0';
				when "01010" => -- BTEQZ
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "010";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '0';
					memoryRead <= '0';
				when "01011" => -- CMP
					aluOp <= "100";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "00";
					regWrite <= '1';
					memoryRead <= '0';
				when "01100" => -- JR
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "100";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '0';
					memoryRead <= '0';
				when "01101" => -- LI
					aluOp <= "111";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '1';
					memoryRead <= '0';
				when "01110" => -- LW
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '0';
					memoryMode <= "10";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '1';
				when "01111" => -- LW_SP
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '0';
					memoryMode <= "10";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '1';
				when "10000" => -- MFIH
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '1';
					memoryRead <= '0';
				when "10001" => -- MFPC
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '1';
					memoryRead <= '0';
				when "10010" => -- MOVE
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '1';
					memoryRead <= '0';
				when "10011" => -- MTIH
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '1';
					memoryRead <= '0';
				when "10100" => -- MTSP
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "11";
					regWrite <= '1';
					memoryRead <= '0';
				when "10101" => -- NOP
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '0';
					memoryRead <= '0';
				when "10110" => -- OR
					aluOp <= "011";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "10111" => -- SLL
					aluOp <= "101";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "11000" => -- SLT
					aluOp <= "001";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "01";
					regWrite <= '1';
					memoryRead <= '0';
				when "11001" => -- SLTI
					aluOp <= "001";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "01";
					regWrite <= '1';
					memoryRead <= '0';
				when "11010" => -- SRA
					aluOp <= "110";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "11011" => -- SUBU
					aluOp <= "001";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '1';
					memoryRead <= '0';
				when "11100" => -- SW
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "01";
					aluResultSrc <= "10";
					regWrite <= '0';
					memoryRead <= '0';
				when "11101" => -- SW_RS
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "01";
					aluResultSrc <= "10";
					regWrite <= '0';
					memoryRead <= '0';
				when "11110" => -- SW_SP
					aluOp <= "000";
					BMuxOp <= '1';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "01";
					aluResultSrc <= "10";
					regWrite <= '0';
					memoryRead <= '0';
				when others => -- NOP
					aluOp <= "111";
					BMuxOp <= '0';
					jumpType <= "000";
					resultSrc <= '1';
					memoryMode <= "00";
					aluResultSrc <= "10";
					regWrite <= '0';
					memoryRead <= '0';
			end case;
		end if;
	end process;
end Behavioral;