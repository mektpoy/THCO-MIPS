library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity MEM2WB is 
    Port ( 
        clk: in STD_LOGIC;
        rst: in STD_LOGIC;
        resultIn : in STD_LOGIC_VECTOR(15 downto 0);
        resultOut : out STD_LOGIC_VECTOR(15 downto 0);
        readDataIn : in STD_LOGIC_VECTOR(15 downto 0);
        readDataOut : out STD_LOGIC_VECTOR(15 downto 0);
        regWbAddrIn : in STD_LOGIC_VECTOR (3 downto 0);
        regWbAddrOut : out STD_LOGIC_VECTOR (3 downto 0);

        --W
        resultSrcIn : in STD_LOGIC;
        resultSrcOut : out STD_LOGIC;
        regWriteClkIn : in STD_LOGIC;
        regWriteClkOut : out STD_LOGIC
    );
end MEM2WB;

architecture Behavioral of MEM2WB is
begin
    process(clk, rst)
    begin
        if(rst = '0') then
            readDataOut <= "0000000000000000";
            resultOut <= "0000000000000000";
            regWbAddrOut <= "0000";
            resultSrcOut <= "0";
            regWriteClkOut <= "0";

        elsif(clk 'event and clk = '1') then
            readDataOut <= readDataIn;
            aluResultOut <= aluResultIn;
            regWbAddrOut <= regWbAddrIn;
            resultSrcOut <= resultSrcIn;
            regWriteClkOut <= regWriteClkIn;
        end if;
    end process;
end Behavioral;